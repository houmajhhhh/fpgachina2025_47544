`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/07/29 14:36:10
// Design Name: 
// Module Name: iic_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module i2c_top (
    input        Clk,
    input        Rst_n,
    input  [7:0] data,
    input        rx_valid,
    
    output       i2c_sclk,
    inout        i2c_sdat,
    output       R_Done,
    output       W_Done,
    output  reg     iic_busy,
    output [7:0] rddata

);

    // �ڲ��ź�����
    
    reg  [7:0]  wrdata;
    reg  [7:0]  device_id_reg;
    reg  [15:0] reg_addr_reg;
    reg  [2:0]  current_state;
    reg  [1:0]  byte_cnt;
    //reg  [7:0]  cmd_buffer [0:2];
    reg         wrreg_req, rdreg_req;
    reg  [15:0] addr;
  //  reg         addr_mode;
   
    
    // ״̬������
    localparam 
        IDLE      = 3'b000,
        CMD_W     = 3'b001,
        CMD_R     = 3'b010,
        CMD_I     = 3'b011;
        //CMD_A     = 3'b100;
    
    reg [2:0] next_state;
    
    // �ֽڼ������߼�
    always @(posedge Clk or negedge Rst_n) begin   //����������  0  ��1��2��0
        if (!Rst_n) begin
            byte_cnt <= 2'b00;
        end else if (rx_valid) begin
            if (byte_cnt == 2'b11)
                byte_cnt <= 2'b00;
            else
                byte_cnt <= byte_cnt + 1'b1;
        end
    end
    
    // ��������洢
//    always @(posedge Clk or negedge Rst_n) begin
//        if (!Rst_n) begin
//            cmd_buffer[0] <= 8'h00;
//            cmd_buffer[1] <= 8'h00;
//            cmd_buffer[2] <= 8'h00;
//        end else if (rx_valid) begin
//            cmd_buffer[byte_cnt] <= data;
//        end
//    end
    
    // ״̬�������߼�
    always @(posedge Clk or negedge Rst_n) begin
        if (!Rst_n) begin
            current_state <= IDLE;
        end else begin
            current_state <= next_state;
        end
    end
    
    // ״̬ת���߼�
    always @(posedge Clk ) begin
        case (current_state)
            IDLE: 
                if ((rx_valid) && (byte_cnt == 2'b00)) begin    //00��01
                    case (data)
                        8'h57: next_state <= CMD_W; // 'W'
                        8'h52: next_state <= CMD_R; // 'R'
                        8'h49: next_state <= CMD_I; // 'I'
                      //  8'h41: next_state = CMD_A; // 'A'
                        default: next_state <= IDLE;
                    endcase
                end else begin
                    next_state = IDLE;
                end
                
            CMD_W: 
                if (rx_valid && byte_cnt == 2'b11)  ///10��00
                    next_state = IDLE;
                else
                    next_state = CMD_W;
                    
            CMD_R: 
                if (rx_valid && byte_cnt == 2'b11)
                    next_state = IDLE;
                else
                    next_state = CMD_R;
                    
            CMD_I: 
                if (rx_valid && byte_cnt == 2'b11)
                    next_state = IDLE;
                else
                    next_state = CMD_I;
                    
//            CMD_A: 
//                if (rx_valid && byte_cnt == 2'b00)
//                    next_state = IDLE;
//                else
//                    next_state = CMD_A;
                    
            default: next_state = IDLE;
        endcase
    end
    
    // �Ĵ�����ַģʽ����
//    always @(posedge Clk or negedge Rst_n) begin
//        if (!Rst_n) begin
//            addr_mode <= 1'b0;
//        end else if (current_state == CMD_A && rx_valid && byte_cnt == 2'b00) begin
//            addr_mode <= data[0]; // ��ַģʽλ
//        end
//    end
    
    // �豸��ַ�Ĵ�������
    always @(posedge Clk or negedge Rst_n) begin
        if (!Rst_n) begin
            device_id_reg <= 8'h00; // Ĭ���豸��ַ
        end else if (current_state == CMD_I && rx_valid && byte_cnt == 2'b01) begin
            device_id_reg <= data;
        end
    end
    
    // �Ĵ�����ַ�Ĵ�������
    always @(posedge Clk or negedge Rst_n) begin
        if (!Rst_n) begin
            reg_addr_reg <= 16'h0000;
        end else if ((current_state == CMD_W||current_state == CMD_R) && rx_valid) begin
            case (byte_cnt)
                2'b01: reg_addr_reg[15:8] <= data;
                2'b10: reg_addr_reg[7:0]  <= data;
                default: ;
            endcase
        end
    end
    
    // I2C������������
    always @(posedge Clk or negedge Rst_n) begin
        if (!Rst_n) begin
            wrreg_req <= 1'b0;
            rdreg_req <= 1'b0;
            addr      <= 16'h0000;
            wrdata    <= 8'h00;
            iic_busy <= 1'b0;
        end else if (current_state == CMD_W && rx_valid && byte_cnt == 2'b11) begin
                wrreg_req <= 1'b1;
              //  addr      <= reg_addr_reg;
                wrdata    <= data;
                iic_busy <=1;
        end else if (current_state == CMD_R && rx_valid && byte_cnt == 2'b11) begin
                rdreg_req <= 1'b1;
                iic_busy <=1;
              //  addr      <= reg_addr_reg;
        end  else if ((iic_busy==1)&&(R_Done==1||W_Done==1)) begin
         wrreg_req <= 1'b0;
         rdreg_req <= 1'b0;   
         iic_busy <= 1'b0;
        end else begin
        wrreg_req <= 1'b0;
        rdreg_req <= 1'b0; 
         end
    end
    
//      always @(posedge Clk or negedge Rst_n) begin
//        if (!Rst_n) begin
//            iic_busy <= 1'b0;
//        end else if ((iic_busy==1)&&(R_Done==1||W_Done==1))
//           iic_busy <= 1'b0;
//        end
        
    // ʵ����I2C������
    i2c_control i2c_control_inst (
        .Clk        (Clk),
        .Rst_n      (Rst_n),
        .wrreg_req  (wrreg_req),
        .rdreg_req  (rdreg_req),
        .addr       (reg_addr_reg),
        .addr_mode  (0),
        .wrdata     (wrdata),
        .rddata     (rddata),
        .device_id  (device_id_reg),
        .R_Done    (R_Done),
        .W_Done    (W_Done),
        .ack        (),
        .i2c_sclk   (i2c_sclk),
        .i2c_sdat   (i2c_sdat)
    );

endmodule