`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/07/24 19:39:10
// Design Name: 
// Module Name: fifo
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module async_fifo #(
    parameter DATA_WIDTH = 8,      // ����λ��
    parameter ADDR_WIDTH = 4       // ��ַλ��2^4=16���
)(
    // д�˿ڣ�дʱ����
    input  wire              wr_clk,     // дʱ��
    input  wire              wr_rst_n,   // д��λ������Ч��
    input  wire              wr_en,      // дʹ��
    input  wire [DATA_WIDTH-1:0] wr_data, // д������
    
    // ���˿ڣ���ʱ����
    input  wire              rd_clk,     // ��ʱ��
    input  wire              rd_rst_n,   // ����λ������Ч��
    input  wire              rd_en,      // ��ʹ��
    output reg  [DATA_WIDTH-1:0] rd_data, // ��������
    
    // ״̬��־
    output wire             full,       // FIFO����־��дʱ����
    output wire             empty       // FIFO�ձ�־����ʱ����
);

    // �ڲ��ź�����
    reg [ADDR_WIDTH:0] wr_ptr_bin;      // дָ�루�����ƣ�
    reg [ADDR_WIDTH:0] rd_ptr_bin;      // ��ָ�루�����ƣ�
    reg [ADDR_WIDTH:0] wr_ptr_gray;     // дָ�루�����룩
    reg [ADDR_WIDTH:0] rd_ptr_gray;     // ��ָ�루�����룩
    
    reg [ADDR_WIDTH:0] rd_ptr_gray_sync1; // ͬ����дʱ����Ķ�ָ�루��һ����
    reg [ADDR_WIDTH:0] rd_ptr_gray_sync2; // ͬ����дʱ����Ķ�ָ�루�ڶ�����
    
    reg [ADDR_WIDTH:0] wr_ptr_gray_sync1; // ͬ������ʱ�����дָ�루��һ����
    reg [ADDR_WIDTH:0] wr_ptr_gray_sync2; // ͬ������ʱ�����дָ�루�ڶ�����
    
    // ˫�˿�RAM�洢����
    reg [DATA_WIDTH-1:0] fifo_mem [0:(1<<ADDR_WIDTH)-1];
    
    // ������ת������
    function [ADDR_WIDTH:0] bin_to_gray(input [ADDR_WIDTH:0] bin);
        bin_to_gray = bin ^ (bin >> 1);
    endfunction
    
    // ������ת������
    function [ADDR_WIDTH:0] gray_to_bin(input [ADDR_WIDTH:0] gray);
        integer i;
        reg [ADDR_WIDTH:0] bin;
        begin
            bin = gray;
            for (i = 1; i <= ADDR_WIDTH; i = i + 1)
                bin = bin ^ (gray >> i);
            gray_to_bin = bin;
        end
    endfunction
    
    // д����
    always @(posedge wr_clk or negedge wr_rst_n) begin
        if (!wr_rst_n) begin
            wr_ptr_bin <= 0;
            wr_ptr_gray <= 0;
        end else if (wr_en && !full) begin
            fifo_mem[wr_ptr_bin[ADDR_WIDTH-1:0]] <= wr_data;
            wr_ptr_bin <= wr_ptr_bin + 1;
            wr_ptr_gray <= bin_to_gray(wr_ptr_bin + 1);
        end
    end
    
    // ������
    always @(posedge rd_clk or negedge rd_rst_n) begin
        if (!rd_rst_n) begin
            rd_ptr_bin <= 0;
            rd_ptr_gray <= 0;
            rd_data <= 0;
        end else if (rd_en && !empty) begin
            rd_data <= fifo_mem[rd_ptr_bin[ADDR_WIDTH-1:0]];
            rd_ptr_bin <= rd_ptr_bin + 1;
            rd_ptr_gray <= bin_to_gray(rd_ptr_bin + 1);
        end
    end
    
    // ��ָ��ͬ����дʱ���������ж���״̬��
    always @(posedge wr_clk or negedge wr_rst_n) begin
        if (!wr_rst_n) begin
            rd_ptr_gray_sync1 <= 0;
            rd_ptr_gray_sync2 <= 0;
        end else begin
            rd_ptr_gray_sync1 <= rd_ptr_gray;
            rd_ptr_gray_sync2 <= rd_ptr_gray_sync1;
        end
    end
    
    // дָ��ͬ������ʱ���������жϿ�״̬��
    always @(posedge rd_clk or negedge rd_rst_n) begin
        if (!rd_rst_n) begin
            wr_ptr_gray_sync1 <= 0;
            wr_ptr_gray_sync2 <= 0;
        end else begin
            wr_ptr_gray_sync1 <= wr_ptr_gray;
            wr_ptr_gray_sync2 <= wr_ptr_gray_sync1;
        end
    end
    
    // ��״̬�жϣ�дʱ����
    assign full = (wr_ptr_gray == {~rd_ptr_gray_sync2[ADDR_WIDTH:ADDR_WIDTH-1], 
                                    rd_ptr_gray_sync2[ADDR_WIDTH-2:0]});
    
    // ��״̬�жϣ���ʱ����
    assign empty = (rd_ptr_gray == wr_ptr_gray_sync2);

endmodule
